`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:18:19 02/26/2019 
// Design Name: 
// Module Name:    top_module 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module top_module(clk, rst, rotate, anode, cathode, mod8Count, inVal, hexVal);

	input wire clk, rst;
	input wire [31:0] inVal;
	wire rotate;
	wire [2:0] mod8Count;
	
	
    );


endmodule
